module ABP_decoder(input a,input b, input c,input clk,input res, output Y, output W );
wire a,b,c,,clk,res;
reg Y,W;  
assign c = 
endmodule
